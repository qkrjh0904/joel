library verilog;
use verilog.vl_types.all;
entity Inen4bit_tb is
end Inen4bit_tb;
