library verilog;
use verilog.vl_types.all;
entity Fourbit_Mul_tb is
end Fourbit_Mul_tb;
