library verilog;
use verilog.vl_types.all;
entity Fourbit_multiplier_tb is
end Fourbit_multiplier_tb;
