library verilog;
use verilog.vl_types.all;
entity InenOen8bit_tb is
end InenOen8bit_tb;
