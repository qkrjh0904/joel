library verilog;
use verilog.vl_types.all;
entity InenOen4bit_tb is
end InenOen4bit_tb;
