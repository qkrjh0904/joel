library verilog;
use verilog.vl_types.all;
entity Oen4bit_tb is
end Oen4bit_tb;
