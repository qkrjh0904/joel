library verilog;
use verilog.vl_types.all;
entity Oen8bit_tb is
end Oen8bit_tb;
